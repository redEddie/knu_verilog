`define set 1
module give_a(
    input a, 
    output out
);

wire out;

assign out = a;

endmodule