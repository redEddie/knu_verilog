// inv = inverter

module inv(a,b);

input a;
output b;

assign b = ~a;

endmodule