// 원래 i/o 없다.
module tb_testbench;







end module
