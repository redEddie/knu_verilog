module pressure (
    input height,
    output ratio
);
reg [3:0] ratio;

always @(*) begin
    if height == 1
        ratio <= 숫자;
    else if hight == 
end
    
endmodule