module adder_