// 정보통신전자공학부 200421379 김철호
// 마이크로 프로세서 설계 기말고사
// Testbench

`timescale 1ns / 1ps
module mut_tb;

	reg clk, rstn, start, load;
	reg [9:0]A, B;
	wire udf, ovf, done;
	wire [9:0]F;

	mut UUT (
		.clk(clk),
		.rstn(rstn),
		.start(start),
		.load(load),
		.A(A),
		.B(B),
		.udf(udf),
		.ovf(ovf),
		.done(done),
		.F(F));

	initial begin 
		clk=0;	rstn=0;start=0; load=0;	
		
		// 기본 연산 테스트
		A=10'b010000_0000;						//    010000_0000	0.1x2^0
		B=10'b010000_0000;						// x 010000_0000	0.1x2^0
		#15 rstn=1;									// --------------------
		#10 load=1;									//    010000_1111	0.01x2^0 => 0.1x2^-1
		#10 start=1 ; load=0;
		#10 start=0;
		
		#60 load=1;
		A=10'b010000_0000;						//    010000_0000	0.1x2^0
		B=10'b010000_1111;						// x 010000_1111	0.1x2^-1
		#10 start=1; load=0;					 	// --------------------
		#10 start=0;									//    010000_1110	0.01x2^-1 => 0.1x2^-2
		
		#60; load=1;
		A=10'b010000_0001;						//    010000_0001	0.1x2^1
		B=10'b010000_0001;						// x 010000_0001  0.1x2^1
		#10 start=1; load=0;					 	// --------------------
		#10 start=0;									//    010000_0001	0.01x2^2 => 0.1x2^1
		
		#60; load=1;
		A=10'b010000_0010;						//    010000_0010	0.1x2^2
		B=10'b010000_0010;						// x 010000_0010  0.1x2^2
		#10 start=1; load=0;					 	// --------------------
		#10 start=0;									//    010000_0011	0.01x2^4 => 0.1x2^3
		
		// 오버 플로우 테스트
		// 양수+양수의 경우 오버 플로우 발생 가능성이 있다.
		#60; load=1;
		A=10'b010000_0101;						//    010000_0101	0.1x2^5
		B=10'b010000_0101;						// x 010000_0101  0.1x2^5
		#10 start=1; load=0;					 	// --------------------
		#10 start=0;									//    010000_1010	0.01x2^10 => 0.1x2^9 => 0.1x2^8 (지수가 8로 오버플로우 발생)
		
		// 언더 플로우 테스트
		// 음수+양수(|양수|<|음수|) 또는 음수+음수의 경우 언더 플로우 발생 가능성이 있다.
		#60; load=1;
		A=10'b010000_1010;						//    010000_1010	0.1x2^-5
		B=10'b010000_1010;						// x 010000_1010  0.1x2^-5
		#10 start=1; load=0;					 	// --------------------
		#10 start=0;									//    010000_1000	0.01x2^-10 => 0.1x2^-11 => 0.1x2^-8 (지수가 -9로 언더플로우 발생)
		
		// 0이 나오는 경우
		#60; load=1;
		A=10'b000000_0011;						//    000000_0011	0.0x2^3
		B=10'b010000_0010;						// x 010000_0010  0.1x2^2
		#10 start=1; load=0;					 	// --------------------
		#10 start=0;									//    000000_0101	0.0x2^5 => 0.0x2^-8  (가수가 0이므로 그냥 제로 처리)
	end
	
	always #5 clk=~clk;
	

endmodule
